
// 3. Behavioural Modeling
module comp1bfull(
    input wire a,
    input wire b,
    output reg c, //As used in an always block need to assign in a reg type
    output reg agb,
    output reg,
);

always @(*) begin // always is used normally in sequential ccts, state machines
    if(a == b) begin
        c = 
    else nota = 1; // else set nota to 1
  
end

endmodule
