module IC7485(
    input wire a,
    input wire b,
    output wire c
);


always @(*) begin
  if (a == b)
end
// can also use
// assign z = (~x & ~y) | (x & y);



endmodule